* Simple LED test circuit
VCC 1 0 DC 5.0
V_IN Q1 0 PULSE(0 5 0ms 0ms 50ms 100ms)
R_OUT Q1 LED_ANODE 50
D1 LED_ANODE LED_CATHODE D_LED
R_LIMIT LED_CATHODE 0 150

.MODEL D_LED D(Is=1e-10 Rs=1 N=1.8 Cjo=10p)

.TRAN 10u 50m
.PRINT TRAN I(D1) V(LED_ANODE) V(LED_CATHODE)
.END
